import "DPI-C" function int factorial(input int i);

program automatic test;
    initial begin
        for (int i=1; i<=10; i++)
            $display("%2d! = %0d", i, factorial(i));
    end
endprogram
